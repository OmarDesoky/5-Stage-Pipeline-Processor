LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY Brach_Forwarding_Unit IS  
PORT (
	--ALU_OUT_EX_MEM,ALU_OUT_2_EX_MEM,MEM_OUT_MEM_WB : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	JMP_SRC,SRC1_EX_MEM,DST_EX_MEM,DST_MEM_WB : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	WB_SIG_EX_MEM, SWAP_SIG_EX_MEM, WB_SIG_MEM_WB,RET_CALL_RTI_READY : IN STD_LOGIC;
	SELECTOR : OUT STD_LOGIC_VECTOR (1 DOWNTO 0)
);    
END ENTITY Brach_Forwarding_Unit;

ARCHITECTURE behavioral_flow OF Brach_Forwarding_Unit IS
BEGIN   

process (SRC1_EX_MEM,DST_EX_MEM,DST_MEM_WB,WB_SIG_EX_MEM, SWAP_SIG_EX_MEM, WB_SIG_MEM_WB , RET_CALL_RTI_READY)
begin
IF (RET_CALL_RTI_READY = '1')
SELECTOR<="11";
ELSIF (JMP_SRC = DST_EX_MEM AND WB_SIG_EX_MEM ='1')THEN
SELECTOR<="01";
ELSIF (JMP_SRC = SRC1_EX_MEM AND WB_SIG_EX_MEM ='1' AND SWAP_SIG_EX_MEM = '1')THEN
SELECTOR<="10";
ELSIF (JMP_SRC = DST_MEM_WB AND WB_SIG_MEM_WB = '1')THEN
SELECTOR<="11";
ELSE 
SELECTOR<="00";
END IF; 
end process;
END behavioral_flow;