LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY Branch_Hazard_Predection_Unit IS  
PORT (
	SRC_CURRENT_OPERATION,DST_ID_EX,DST_EX_MEM,INSTRCTION_10_8_DECODE_STAGE,INSTRUCTION_7_5_DECODE_STAGE,INSTRUCTION_4_2_DECODE_STAGE,SRC1_ID_EX,
	SRC2_ID_EX : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	ENABLE,WB_SIG_DECODE_STAGE,WB_SIG_ID_EX,SWAP_SIG_DECODE_STAGE,SWAP_SIG_ID_EX,MEM_READ_SIG_DECODE_STAGE,MEM_READ_ID_EX,MEM_READ_EX_MEM,WB_SIG_EX_MEM : IN STD_LOGIC;
	STALL_SIGNAL : OUT STD_LOGIC
);    
END ENTITY Branch_Hazard_Predection_Unit;

ARCHITECTURE behavioral_flow OF Branch_Hazard_Predection_Unit IS
BEGIN   

process (SRC_CURRENT_OPERATION,DST_ID_EX,DST_EX_MEM,INSTRCTION_10_8_DECODE_STAGE,INSTRUCTION_7_5_DECODE_STAGE,INSTRUCTION_4_2_DECODE_STAGE,SRC1_ID_EX,
	SRC2_ID_EX,ENABLE,WB_SIG_DECODE_STAGE,WB_SIG_ID_EX,SWAP_SIG_DECODE_STAGE,SWAP_SIG_ID_EX,MEM_READ_SIG_DECODE_STAGE,MEM_READ_ID_EX,MEM_READ_EX_MEM,WB_SIG_EX_MEM)
begin
IF (ENABLE = '1')
THEN
	STALL_SIGNAL <= '0';

	-- CASE SWAP IN THE DECODE STAGE
	IF (WB_SIG_DECODE_STAGE = '1' AND (SRC_CURRENT_OPERATION = INSTRUCTION_7_5_DECODE_STAGE OR SRC_CURRENT_OPERATION = INSTRUCTION_4_2_DECODE_STAGE )AND SWAP_SIG_DECODE_STAGE = '1')
	THEN 
		STALL_SIGNAL <= '1';
	-- CASE SWAP IN THE EXECUTE STAGE
	ELSIF (WB_SIG_ID_EX = '1' AND (SRC_CURRENT_OPERATION = SRC1_ID_EX OR SRC_CURRENT_OPERATION = SRC2_ID_EX )AND SWAP_SIG_ID_EX = '1')
	THEN 
		STALL_SIGNAL <= '1';

	-- CASE LDD IN DECODE STAGE
	ELSIF (WB_SIG_DECODE_STAGE = '1' AND MEM_READ_SIG_DECODE_STAGE = '1' AND SRC_CURRENT_OPERATION = DST_ID_EX)
	THEN 
		STALL_SIGNAL <= '1';
	-- CASE LDD IN EXECUTE STAGE
	ELSIF (WB_SIG_ID_EX = '1' AND MEM_READ_ID_EX = '1' AND SRC_CURRENT_OPERATION = DST_ID_EX)
	THEN 
		STALL_SIGNAL <= '1';
	-- CASE LDD IN MEMORY STAGE
	ELSIF (WB_SIG_EX_MEM = '1' AND MEM_READ_EX_MEM = '1' AND SRC_CURRENT_OPERATION = DST_EX_MEM)
	THEN 
		STALL_SIGNAL <= '1';
	-- CASE LDM & 1_OPERAND IN 2ND CYCLE IN DECODE
	ELSIF (WB_SIG_DECODE_STAGE = '1' AND (SRC_CURRENT_OPERATION = DST_ID_EX OR SRC_CURRENT_OPERATION = INSTRCTION_10_8_DECODE_STAGE))
	THEN 
		STALL_SIGNAL <= '1';
	-- CASE LDM & 1_OPERAND IN EXECUTION
	ELSIF (WB_SIG_ID_EX = '1' AND SRC_CURRENT_OPERATION = DST_ID_EX)
	THEN 
		STALL_SIGNAL <= '1';
	END IF;
ELSE
STALL_SIGNAL <= '0';
END IF;
end process;
END behavioral_flow;